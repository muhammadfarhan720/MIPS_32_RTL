
module AND(e,f,g);

input e,f; 
output  g; 


 
 assign g= e & f ;
 

endmodule