
module AND(e,f,g);

input e,f; 
output reg g; 

always @(*)
 
 g= e & f ;

endmodule